
module SCJIO (
	tms,
	tdi,
	tdo,
	tck);	

	input		tms;
	input		tdi;
	output		tdo;
	input		tck;
endmodule
