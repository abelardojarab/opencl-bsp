package hssi_eth_pkg;
parameter NUM_LN = 16;    
endpackage
