// SCJIO.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module SCJIO (
		input  wire  tms, // jtag.tms
		input  wire  tdi, //     .tdi
		output wire  tdo, //     .tdo
		input  wire  tck  //  tck.clk
	);

	altera_soft_core_jtag_io #(
		.ENABLE_JTAG_IO_SELECTION (0)
	) soft_core_jtag_io_0 (
		.tms         (tms),  // jtag.tms
		.tdi         (tdi),  //     .tdi
		.tdo         (tdo),  //     .tdo
		.tck         (tck),  //  tck.clk
		.select_this (1'b0)  // (terminated)
	);

endmodule
