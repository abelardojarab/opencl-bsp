module global_routing
(
   input s,
   input clk,
   output g
);

assign g = s;

endmodule
