// ***************************************************************************
// Copyright (c) 2013-2017, Intel Corporation All Rights Reserved.
// The source code contained or described herein and all  documents related to
// the  source  code  ("Material")  are  owned by  Intel  Corporation  or  its
// suppliers  or  licensors.    Title  to  the  Material  remains  with  Intel
// Corporation or  its suppliers  and licensors.  The Material  contains trade
// secrets and  proprietary  and  confidential  information  of  Intel or  its
// suppliers and licensors.  The Material is protected  by worldwide copyright
// and trade secret laws and treaty provisions. No part of the Material may be
// copied,    reproduced,    modified,    published,     uploaded,     posted,
// transmitted,  distributed,  or  disclosed  in any way without Intel's prior
// express written permission.
// ***************************************************************************

`ifndef SYS_CFG_PKG_SV                                          
    `define SYS_CFG_PKG_SV      
//  `define CCIP_DEBUG              // Add ccip_debug_module
    `define VENDOR_ALTERA           // Use Altera FPGA
    `define TOOL_QUARTUS            // Use Altera Quartus Tools     
`endif
 

